module InstructionMemory(
	input logic clk,
	input logic [7:0] Address,
	input logic rst,
	output logic [31:0] ReadData
);

	logic [31:0] regData [511:0];

	logic error_addr;


	// TODO: Bit width of the pc addressing
	logic [7:0] direct_addressing;
	assign direct_addressing = Address >> 2;

	assign error_addr = |(Address % 4);

	assign ReadData = regData[direct_addressing];
	

	// //SW$1,0($2)
	// assign regData[0]=32'b10101100010000010000000000000000;
	// //LW$5,0($4)
	// assign regData[1]=32'b10001100100001010000000000000000;
	// //BEQ$5,$1,1
	// assign regData[2]=32'b00010000101000010000000000000001;
	// //JMP1
	// assign regData[3]=32'b00001000000000000000000000000001;

	// //SW $10,0($3)////
	// assign regData[4]=32'b10101100011010100000000000000000;
	// //SW$20,0($1)
	// assign regData[5]=32'b10101110100000010000000000000000;
	// //LW$5,0($21)
	// assign regData[6]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)	
	// assign regData[7]=32'b10101110100000000000000000000000;	
	// //BEQ$5,$1,1
	// assign regData[8]=32'b00010000101000010000000000000001;
	// //JUMP 5
	// assign regData[9]=32'b00001000000000000000000000000101;

	// //LW$11,0($3)
	// assign regData[10]=32'b10101100011010110000000000000000;
	// //SW$20,0($1)
	// assign regData[11]=32'b10101110100000010000000000000000;
	// //LW$5,0($21)
	// assign regData[12]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[13]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[14]=32'b00010000101000010000000000000001;
	// //JUMP11
	// assign regData[15]=32'b00001000000000000000000000001011;

	// //LW$12,0($3)
	// assign regData[16]=32'b10101100011011000000000000000000;
	// //SW$20,0($1)
	// assign regData[17]=32'b10101110100000010000000000000000;	
	// //LW$5,0($21)
	// assign regData[18]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[19]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[20]=32'b00010000101000010000000000000001;
	// //JUMP18
	// assign regData[21]=32'b00001000000000000000000000010001;

	// //LW$13,0($3)   
	// assign regData[22]=32'b10101100011011010000000000000000;
	// //SW$20,0($1)
	// assign regData[23]=32'b10101110100000010000000000000000;	
	// //LW$5,0($21)
	// assign regData[24]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[25]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[26]=32'b00010000101000010000000000000001;
	// //JUMP
	// assign regData[27]=32'b00001000000000000000000000010111;


	// //LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
	// assign regData[28]=32'b10101100011011100000000000000000;
	// //SW$20,0($1)
	// assign regData[29]=32'b10101110100000010000000000000000;	
	// //LW$5,0($21)
	// assign regData[30]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[31]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[32]=32'b00010000101000010000000000000001;
	// //JUMP
	// assign regData[33]=32'b00001000000000000000000000011101;

	// //LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
	// assign regData[34]=32'b10101100011011110000000000000000;
	// //SW$20,0($1)
	// assign regData[35]=32'b10101110100000010000000000000000;	
	// //LW$5,0($21)
	// assign regData[36]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[37]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[38]=32'b00010000101000010000000000000001;
	// //JUMP
	// assign regData[39]=32'b00001000000000000000000000100011;


	// //LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
	// assign regData[40]=32'b10101100011100000000000000000000;
	// //SW$20,0($1)
	// assign regData[41]=32'b10101110100000010000000000000000;	
	// //LW$5,0($21)
	// assign regData[42]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[43]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[44]=32'b00010000101000010000000000000001;
	// //JUMP
	// assign regData[45]=32'b00001000000000000000000000101001;

	// //LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
	// assign regData[46]=32'b10101100011100010000000000000000;
	// //SW$20,0($1)
	// assign regData[47]=32'b10101110100000010000000000000000;	
	// //LW$5,0($21)
	// assign regData[48]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[49]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[50]=32'b00010000101000010000000000000001;
	// //JUMP
	// assign regData[51]=32'b00001000000000000000000000101111;

	// //LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
	// assign regData[52]=32'b10101100011100100000000000000000;
	// //SW$20,0($1)
	// assign regData[53]=32'b10101110100000010000000000000000;	
	// //LW$5,0($21)
	// assign regData[54]=32'b10001110101001010000000000000000;
	// //SW$20,0($0)
	// assign regData[55]=32'b10101110100000000000000000000000;
	// //BEQ$5,$1,1
	// assign regData[56]=32'b00010000101000010000000000000001;
	// //JUMP
	// assign regData[57]=32'b00001000000000000000000000110101;
	// //STAY 
	// assign regData[58]=32'b00001000000000000000000000111010;




endmodule
