module InstructionMemory(
	input clk,
	input [7:0] Address,
	input rst,
	output logic [31:0] ReadData
);

	logic [31:0] regData [511:0];
	
	assign ReadData = regData[Address];
	
	always_ff @ (posedge clk) begin
		if (rst) begin
		 	for(int j = 0; j<512; j= j +1) begin
				regData[j] = 0;
			end
			


				//SW$1,0($2)
				regData[0]=32'b10101100010000010000000000000000;
				//LW$5,0($4)
				regData[1]=32'b10001100100001010000000000000000;
				//BEQ$5,$1,1
				regData[2]=32'b00010000101000010000000000000001;
				//JMP1
				regData[3]=32'b00001000000000000000000000000001;

				//SW $10,0($3)////
				regData[4]=32'b10101100011010100000000000000000;
				//SW$20,0($1)
				regData[5]=32'b10101110100000010000000000000000;
				//LW$5,0($21)
				regData[6]=32'b10001110101001010000000000000000;
				//SW$20,0($0)	
				regData[7]=32'b10101110100000000000000000000000;	
				//BEQ$5,$1,1
				regData[8]=32'b00010000101000010000000000000001;
				//JUMP 5
				regData[9]=32'b00001000000000000000000000000101;

				//LW$11,0($3)
				regData[10]=32'b10101100011010110000000000000000;
				//SW$20,0($1)
				regData[11]=32'b10101110100000010000000000000000;
				//LW$5,0($21)
				regData[12]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[13]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[14]=32'b00010000101000010000000000000001;
				//JUMP11
				regData[15]=32'b00001000000000000000000000001011;

				//LW$12,0($3)
				regData[16]=32'b10101100011011000000000000000000;
				//SW$20,0($1)
				regData[17]=32'b10101110100000010000000000000000;	
				//LW$5,0($21)
				regData[18]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[19]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[20]=32'b00010000101000010000000000000001;
				//JUMP18
				regData[21]=32'b00001000000000000000000000010001;

				//LW$13,0($3)   
				regData[22]=32'b10101100011011010000000000000000;
				//SW$20,0($1)
				regData[23]=32'b10101110100000010000000000000000;	
				//LW$5,0($21)
				regData[24]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[25]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[26]=32'b00010000101000010000000000000001;
				//JUMP
				regData[27]=32'b00001000000000000000000000010111;


				//LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
				regData[28]=32'b10101100011011100000000000000000;
				//SW$20,0($1)
				regData[29]=32'b10101110100000010000000000000000;	
				//LW$5,0($21)
				regData[30]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[31]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[32]=32'b00010000101000010000000000000001;
				//JUMP
				regData[33]=32'b00001000000000000000000000011101;

				//LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
				regData[34]=32'b10101100011011110000000000000000;
				//SW$20,0($1)
				regData[35]=32'b10101110100000010000000000000000;	
				//LW$5,0($21)
				regData[36]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[37]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[38]=32'b00010000101000010000000000000001;
				//JUMP
				regData[39]=32'b00001000000000000000000000100011;


				//LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
				regData[40]=32'b10101100011100000000000000000000;
				//SW$20,0($1)
				regData[41]=32'b10101110100000010000000000000000;	
				//LW$5,0($21)
				regData[42]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[43]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[44]=32'b00010000101000010000000000000001;
				//JUMP
				regData[45]=32'b00001000000000000000000000101001;

				//LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
				regData[46]=32'b10101100011100010000000000000000;
				//SW$20,0($1)
				regData[47]=32'b10101110100000010000000000000000;	
				//LW$5,0($21)
				regData[48]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[49]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[50]=32'b00010000101000010000000000000001;
				//JUMP
				regData[51]=32'b00001000000000000000000000101111;

				//LW$13,0($3)   100011ssssstttttiiiiiiiiiiiiiiii
				regData[52]=32'b10101100011100100000000000000000;
				//SW$20,0($1)
				regData[53]=32'b10101110100000010000000000000000;	
				//LW$5,0($21)
				regData[54]=32'b10001110101001010000000000000000;
				//SW$20,0($0)
				regData[55]=32'b10101110100000000000000000000000;
				//BEQ$5,$1,1
				regData[56]=32'b00010000101000010000000000000001;
				//JUMP
				regData[57]=32'b00001000000000000000000000110101;

				//STAY 
				regData[58]=32'b00001000000000000000000000111010;






			end
	end
	
//	always @ (posedge clk)begin
//		ReadData <= regData[Address];
//	end

endmodule
